QuadTest_12chFF_64B66B.vhd